module memStage(
	input clk,
	input [31:0] alu_result,
	input [31:0] datainput,
	input [4:0] rd,
	input [2:0] flagsMEM,
	input [1:0] flagsWB,
	output [1:0] flagsWB_out,
	output [31:0] mem_data,
	output [31:0] direction,
	output [4:0] rd_out
);

	

	
	assign flagsWB_out = flagsWB;
	assign direction = alu_result;
	assign rd_out = rd;

endmodule